* C:\Users\kesav\eSim-Workspace\finaltry\finaltry.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/22/20 10:36:15

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  sample Net-_M2-Pad2_ input input eSim_MOS_P		
M1  input Net-_M1-Pad2_ sample sample eSim_MOS_N		
X1  Net-_M1-Pad2_ Net-_M2-Pad2_ INVCMOS		
v1  input GND sine		
v2  Net-_M1-Pad2_ GND pulse		
C1  sample GND .1u		
U2  sample plot_v1		
U1  input plot_v1		
R3  ? GND 2k		

.end
